module rom_lut_sin (
    input clk, rst_n,
    input [8:0] addr_i,
    output reg signed [15:0] value_o
);

always@(posedge clk or negedge rst_n)
    if(!rst_n)
        value_o <= 'd0 ;  
    else  begin
      case(addr_i) 
9'd0:value_o <=    16'd0;
9'd1:value_o <=    16'd402;
9'd2:value_o <=    16'd804;
9'd3:value_o <=    16'd1206;
9'd4:value_o <=    16'd1608;
9'd5:value_o <=    16'd2009;
9'd6:value_o <=    16'd2411;
9'd7:value_o <=    16'd2811;
9'd8:value_o <=    16'd3212;
9'd9:value_o <=    16'd3612;
9'd10:value_o <=    16'd4011;
9'd11:value_o <=    16'd4410;
9'd12:value_o <=    16'd4808;
9'd13:value_o <=    16'd5205;
9'd14:value_o <=    16'd5602;
9'd15:value_o <=    16'd5998;
9'd16:value_o <=    16'd6393;
9'd17:value_o <=    16'd6787;
9'd18:value_o <=    16'd7179;
9'd19:value_o <=    16'd7571;
9'd20:value_o <=    16'd7962;
9'd21:value_o <=    16'd8351;
9'd22:value_o <=    16'd8740;
9'd23:value_o <=    16'd9126;
9'd24:value_o <=    16'd9512;
9'd25:value_o <=    16'd9896;
9'd26:value_o <=    16'd10279;
9'd27:value_o <=    16'd10660;
9'd28:value_o <=    16'd11039;
9'd29:value_o <=    16'd11417;
9'd30:value_o <=    16'd11793;
9'd31:value_o <=    16'd12167;
9'd32:value_o <=    16'd12540;
9'd33:value_o <=    16'd12910;
9'd34:value_o <=    16'd13279;
9'd35:value_o <=    16'd13645;
9'd36:value_o <=    16'd14010;
9'd37:value_o <=    16'd14372;
9'd38:value_o <=    16'd14733;
9'd39:value_o <=    16'd15091;
9'd40:value_o <=    16'd15446;
9'd41:value_o <=    16'd15800;
9'd42:value_o <=    16'd16151;
9'd43:value_o <=    16'd16500;
9'd44:value_o <=    16'd16846;
9'd45:value_o <=    16'd17189;
9'd46:value_o <=    16'd17531;
9'd47:value_o <=    16'd17869;
9'd48:value_o <=    16'd18205;
9'd49:value_o <=    16'd18538;
9'd50:value_o <=    16'd18868;
9'd51:value_o <=    16'd19195;
9'd52:value_o <=    16'd19520;
9'd53:value_o <=    16'd19841;
9'd54:value_o <=    16'd20160;
9'd55:value_o <=    16'd20475;
9'd56:value_o <=    16'd20787;
9'd57:value_o <=    16'd21097;
9'd58:value_o <=    16'd21403;
9'd59:value_o <=    16'd21706;
9'd60:value_o <=    16'd22005;
9'd61:value_o <=    16'd22302;
9'd62:value_o <=    16'd22595;
9'd63:value_o <=    16'd22884;
9'd64:value_o <=    16'd23170;
9'd65:value_o <=    16'd23453;
9'd66:value_o <=    16'd23732;
9'd67:value_o <=    16'd24007;
9'd68:value_o <=    16'd24279;
9'd69:value_o <=    16'd24547;
9'd70:value_o <=    16'd24812;
9'd71:value_o <=    16'd25073;
9'd72:value_o <=    16'd25330;
9'd73:value_o <=    16'd25583;
9'd74:value_o <=    16'd25832;
9'd75:value_o <=    16'd26078;
9'd76:value_o <=    16'd26319;
9'd77:value_o <=    16'd26557;
9'd78:value_o <=    16'd26790;
9'd79:value_o <=    16'd27020;
9'd80:value_o <=    16'd27245;
9'd81:value_o <=    16'd27467;
9'd82:value_o <=    16'd27684;
9'd83:value_o <=    16'd27897;
9'd84:value_o <=    16'd28106;
9'd85:value_o <=    16'd28310;
9'd86:value_o <=    16'd28511;
9'd87:value_o <=    16'd28707;
9'd88:value_o <=    16'd28898;
9'd89:value_o <=    16'd29086;
9'd90:value_o <=    16'd29269;
9'd91:value_o <=    16'd29447;
9'd92:value_o <=    16'd29621;
9'd93:value_o <=    16'd29791;
9'd94:value_o <=    16'd29956;
9'd95:value_o <=    16'd30117;
9'd96:value_o <=    16'd30273;
9'd97:value_o <=    16'd30425;
9'd98:value_o <=    16'd30572;
9'd99:value_o <=    16'd30714;
9'd100:value_o <=    16'd30852;
9'd101:value_o <=    16'd30985;
9'd102:value_o <=    16'd31114;
9'd103:value_o <=    16'd31237;
9'd104:value_o <=    16'd31357;
9'd105:value_o <=    16'd31471;
9'd106:value_o <=    16'd31581;
9'd107:value_o <=    16'd31685;
9'd108:value_o <=    16'd31785;
9'd109:value_o <=    16'd31881;
9'd110:value_o <=    16'd31971;
9'd111:value_o <=    16'd32057;
9'd112:value_o <=    16'd32138;
9'd113:value_o <=    16'd32214;
9'd114:value_o <=    16'd32285;
9'd115:value_o <=    16'd32351;
9'd116:value_o <=    16'd32413;
9'd117:value_o <=    16'd32469;
9'd118:value_o <=    16'd32521;
9'd119:value_o <=    16'd32568;
9'd120:value_o <=    16'd32610;
9'd121:value_o <=    16'd32647;
9'd122:value_o <=    16'd32679;
9'd123:value_o <=    16'd32706;
9'd124:value_o <=    16'd32728;
9'd125:value_o <=    16'd32745;
9'd126:value_o <=    16'd32758;
9'd127:value_o <=    16'd32765;
9'd128:value_o <=    16'd32768;
9'd129:value_o <=    16'd32765;
9'd130:value_o <=    16'd32758;
9'd131:value_o <=    16'd32745;
9'd132:value_o <=    16'd32728;
9'd133:value_o <=    16'd32706;
9'd134:value_o <=    16'd32679;
9'd135:value_o <=    16'd32647;
9'd136:value_o <=    16'd32610;
9'd137:value_o <=    16'd32568;
9'd138:value_o <=    16'd32521;
9'd139:value_o <=    16'd32469;
9'd140:value_o <=    16'd32413;
9'd141:value_o <=    16'd32351;
9'd142:value_o <=    16'd32285;
9'd143:value_o <=    16'd32214;
9'd144:value_o <=    16'd32138;
9'd145:value_o <=    16'd32057;
9'd146:value_o <=    16'd31971;
9'd147:value_o <=    16'd31881;
9'd148:value_o <=    16'd31785;
9'd149:value_o <=    16'd31685;
9'd150:value_o <=    16'd31581;
9'd151:value_o <=    16'd31471;
9'd152:value_o <=    16'd31357;
9'd153:value_o <=    16'd31237;
9'd154:value_o <=    16'd31114;
9'd155:value_o <=    16'd30985;
9'd156:value_o <=    16'd30852;
9'd157:value_o <=    16'd30714;
9'd158:value_o <=    16'd30572;
9'd159:value_o <=    16'd30425;
9'd160:value_o <=    16'd30273;
9'd161:value_o <=    16'd30117;
9'd162:value_o <=    16'd29956;
9'd163:value_o <=    16'd29791;
9'd164:value_o <=    16'd29621;
9'd165:value_o <=    16'd29447;
9'd166:value_o <=    16'd29269;
9'd167:value_o <=    16'd29086;
9'd168:value_o <=    16'd28898;
9'd169:value_o <=    16'd28707;
9'd170:value_o <=    16'd28511;
9'd171:value_o <=    16'd28310;
9'd172:value_o <=    16'd28106;
9'd173:value_o <=    16'd27897;
9'd174:value_o <=    16'd27684;
9'd175:value_o <=    16'd27467;
9'd176:value_o <=    16'd27245;
9'd177:value_o <=    16'd27020;
9'd178:value_o <=    16'd26790;
9'd179:value_o <=    16'd26557;
9'd180:value_o <=    16'd26319;
9'd181:value_o <=    16'd26078;
9'd182:value_o <=    16'd25832;
9'd183:value_o <=    16'd25583;
9'd184:value_o <=    16'd25330;
9'd185:value_o <=    16'd25073;
9'd186:value_o <=    16'd24812;
9'd187:value_o <=    16'd24547;
9'd188:value_o <=    16'd24279;
9'd189:value_o <=    16'd24007;
9'd190:value_o <=    16'd23732;
9'd191:value_o <=    16'd23453;
9'd192:value_o <=    16'd23170;
9'd193:value_o <=    16'd22884;
9'd194:value_o <=    16'd22595;
9'd195:value_o <=    16'd22302;
9'd196:value_o <=    16'd22005;
9'd197:value_o <=    16'd21706;
9'd198:value_o <=    16'd21403;
9'd199:value_o <=    16'd21097;
9'd200:value_o <=    16'd20787;
9'd201:value_o <=    16'd20475;
9'd202:value_o <=    16'd20160;
9'd203:value_o <=    16'd19841;
9'd204:value_o <=    16'd19520;
9'd205:value_o <=    16'd19195;
9'd206:value_o <=    16'd18868;
9'd207:value_o <=    16'd18538;
9'd208:value_o <=    16'd18205;
9'd209:value_o <=    16'd17869;
9'd210:value_o <=    16'd17531;
9'd211:value_o <=    16'd17189;
9'd212:value_o <=    16'd16846;
9'd213:value_o <=    16'd16500;
9'd214:value_o <=    16'd16151;
9'd215:value_o <=    16'd15800;
9'd216:value_o <=    16'd15446;
9'd217:value_o <=    16'd15091;
9'd218:value_o <=    16'd14733;
9'd219:value_o <=    16'd14372;
9'd220:value_o <=    16'd14010;
9'd221:value_o <=    16'd13645;
9'd222:value_o <=    16'd13279;
9'd223:value_o <=    16'd12910;
9'd224:value_o <=    16'd12540;
9'd225:value_o <=    16'd12167;
9'd226:value_o <=    16'd11793;
9'd227:value_o <=    16'd11417;
9'd228:value_o <=    16'd11039;
9'd229:value_o <=    16'd10660;
9'd230:value_o <=    16'd10279;
9'd231:value_o <=    16'd9896;
9'd232:value_o <=    16'd9512;
9'd233:value_o <=    16'd9126;
9'd234:value_o <=    16'd8740;
9'd235:value_o <=    16'd8351;
9'd236:value_o <=    16'd7962;
9'd237:value_o <=    16'd7571;
9'd238:value_o <=    16'd7179;
9'd239:value_o <=    16'd6787;
9'd240:value_o <=    16'd6393;
9'd241:value_o <=    16'd5998;
9'd242:value_o <=    16'd5602;
9'd243:value_o <=    16'd5205;
9'd244:value_o <=    16'd4808;
9'd245:value_o <=    16'd4410;
9'd246:value_o <=    16'd4011;
9'd247:value_o <=    16'd3612;
9'd248:value_o <=    16'd3212;
9'd249:value_o <=    16'd2811;
9'd250:value_o <=    16'd2411;
9'd251:value_o <=    16'd2009;
9'd252:value_o <=    16'd1608;
9'd253:value_o <=    16'd1206;
9'd254:value_o <=    16'd804;
9'd255:value_o <=    16'd402;
9'd256:value_o <=    16'd0;
9'd257:value_o <=    16'd65133;
9'd258:value_o <=    16'd64731;
9'd259:value_o <=    16'd64329;
9'd260:value_o <=    16'd63927;
9'd261:value_o <=    16'd63526;
9'd262:value_o <=    16'd63124;
9'd263:value_o <=    16'd62724;
9'd264:value_o <=    16'd62323;
9'd265:value_o <=    16'd61923;
9'd266:value_o <=    16'd61524;
9'd267:value_o <=    16'd61125;
9'd268:value_o <=    16'd60727;
9'd269:value_o <=    16'd60330;
9'd270:value_o <=    16'd59933;
9'd271:value_o <=    16'd59537;
9'd272:value_o <=    16'd59142;
9'd273:value_o <=    16'd58748;
9'd274:value_o <=    16'd58356;
9'd275:value_o <=    16'd57964;
9'd276:value_o <=    16'd57573;
9'd277:value_o <=    16'd57184;
9'd278:value_o <=    16'd56795;
9'd279:value_o <=    16'd56409;
9'd280:value_o <=    16'd56023;
9'd281:value_o <=    16'd55639;
9'd282:value_o <=    16'd55256;
9'd283:value_o <=    16'd54875;
9'd284:value_o <=    16'd54496;
9'd285:value_o <=    16'd54118;
9'd286:value_o <=    16'd53742;
9'd287:value_o <=    16'd53368;
9'd288:value_o <=    16'd52995;
9'd289:value_o <=    16'd52625;
9'd290:value_o <=    16'd52256;
9'd291:value_o <=    16'd51890;
9'd292:value_o <=    16'd51525;
9'd293:value_o <=    16'd51163;
9'd294:value_o <=    16'd50802;
9'd295:value_o <=    16'd50444;
9'd296:value_o <=    16'd50089;
9'd297:value_o <=    16'd49735;
9'd298:value_o <=    16'd49384;
9'd299:value_o <=    16'd49035;
9'd300:value_o <=    16'd48689;
9'd301:value_o <=    16'd48346;
9'd302:value_o <=    16'd48004;
9'd303:value_o <=    16'd47666;
9'd304:value_o <=    16'd47330;
9'd305:value_o <=    16'd46997;
9'd306:value_o <=    16'd46667;
9'd307:value_o <=    16'd46340;
9'd308:value_o <=    16'd46015;
9'd309:value_o <=    16'd45694;
9'd310:value_o <=    16'd45375;
9'd311:value_o <=    16'd45060;
9'd312:value_o <=    16'd44748;
9'd313:value_o <=    16'd44438;
9'd314:value_o <=    16'd44132;
9'd315:value_o <=    16'd43829;
9'd316:value_o <=    16'd43530;
9'd317:value_o <=    16'd43233;
9'd318:value_o <=    16'd42940;
9'd319:value_o <=    16'd42651;
9'd320:value_o <=    16'd42365;
9'd321:value_o <=    16'd42082;
9'd322:value_o <=    16'd41803;
9'd323:value_o <=    16'd41528;
9'd324:value_o <=    16'd41256;
9'd325:value_o <=    16'd40988;
9'd326:value_o <=    16'd40723;
9'd327:value_o <=    16'd40462;
9'd328:value_o <=    16'd40205;
9'd329:value_o <=    16'd39952;
9'd330:value_o <=    16'd39703;
9'd331:value_o <=    16'd39457;
9'd332:value_o <=    16'd39216;
9'd333:value_o <=    16'd38978;
9'd334:value_o <=    16'd38745;
9'd335:value_o <=    16'd38515;
9'd336:value_o <=    16'd38290;
9'd337:value_o <=    16'd38068;
9'd338:value_o <=    16'd37851;
9'd339:value_o <=    16'd37638;
9'd340:value_o <=    16'd37429;
9'd341:value_o <=    16'd37225;
9'd342:value_o <=    16'd37024;
9'd343:value_o <=    16'd36828;
9'd344:value_o <=    16'd36637;
9'd345:value_o <=    16'd36449;
9'd346:value_o <=    16'd36266;
9'd347:value_o <=    16'd36088;
9'd348:value_o <=    16'd35914;
9'd349:value_o <=    16'd35744;
9'd350:value_o <=    16'd35579;
9'd351:value_o <=    16'd35418;
9'd352:value_o <=    16'd35262;
9'd353:value_o <=    16'd35110;
9'd354:value_o <=    16'd34963;
9'd355:value_o <=    16'd34821;
9'd356:value_o <=    16'd34683;
9'd357:value_o <=    16'd34550;
9'd358:value_o <=    16'd34421;
9'd359:value_o <=    16'd34298;
9'd360:value_o <=    16'd34178;
9'd361:value_o <=    16'd34064;
9'd362:value_o <=    16'd33954;
9'd363:value_o <=    16'd33850;
9'd364:value_o <=    16'd33750;
9'd365:value_o <=    16'd33654;
9'd366:value_o <=    16'd33564;
9'd367:value_o <=    16'd33478;
9'd368:value_o <=    16'd33397;
9'd369:value_o <=    16'd33321;
9'd370:value_o <=    16'd33250;
9'd371:value_o <=    16'd33184;
9'd372:value_o <=    16'd33122;
9'd373:value_o <=    16'd33066;
9'd374:value_o <=    16'd33014;
9'd375:value_o <=    16'd32967;
9'd376:value_o <=    16'd32925;
9'd377:value_o <=    16'd32888;
9'd378:value_o <=    16'd32856;
9'd379:value_o <=    16'd32829;
9'd380:value_o <=    16'd32807;
9'd381:value_o <=    16'd32790;
9'd382:value_o <=    16'd32777;
9'd383:value_o <=    16'd32770;
9'd384:value_o <=    16'd32768;
9'd385:value_o <=    16'd32770;
9'd386:value_o <=    16'd32777;
9'd387:value_o <=    16'd32790;
9'd388:value_o <=    16'd32807;
9'd389:value_o <=    16'd32829;
9'd390:value_o <=    16'd32856;
9'd391:value_o <=    16'd32888;
9'd392:value_o <=    16'd32925;
9'd393:value_o <=    16'd32967;
9'd394:value_o <=    16'd33014;
9'd395:value_o <=    16'd33066;
9'd396:value_o <=    16'd33122;
9'd397:value_o <=    16'd33184;
9'd398:value_o <=    16'd33250;
9'd399:value_o <=    16'd33321;
9'd400:value_o <=    16'd33397;
9'd401:value_o <=    16'd33478;
9'd402:value_o <=    16'd33564;
9'd403:value_o <=    16'd33654;
9'd404:value_o <=    16'd33750;
9'd405:value_o <=    16'd33850;
9'd406:value_o <=    16'd33954;
9'd407:value_o <=    16'd34064;
9'd408:value_o <=    16'd34178;
9'd409:value_o <=    16'd34298;
9'd410:value_o <=    16'd34421;
9'd411:value_o <=    16'd34550;
9'd412:value_o <=    16'd34683;
9'd413:value_o <=    16'd34821;
9'd414:value_o <=    16'd34963;
9'd415:value_o <=    16'd35110;
9'd416:value_o <=    16'd35262;
9'd417:value_o <=    16'd35418;
9'd418:value_o <=    16'd35579;
9'd419:value_o <=    16'd35744;
9'd420:value_o <=    16'd35914;
9'd421:value_o <=    16'd36088;
9'd422:value_o <=    16'd36266;
9'd423:value_o <=    16'd36449;
9'd424:value_o <=    16'd36637;
9'd425:value_o <=    16'd36828;
9'd426:value_o <=    16'd37024;
9'd427:value_o <=    16'd37225;
9'd428:value_o <=    16'd37429;
9'd429:value_o <=    16'd37638;
9'd430:value_o <=    16'd37851;
9'd431:value_o <=    16'd38068;
9'd432:value_o <=    16'd38290;
9'd433:value_o <=    16'd38515;
9'd434:value_o <=    16'd38745;
9'd435:value_o <=    16'd38978;
9'd436:value_o <=    16'd39216;
9'd437:value_o <=    16'd39457;
9'd438:value_o <=    16'd39703;
9'd439:value_o <=    16'd39952;
9'd440:value_o <=    16'd40205;
9'd441:value_o <=    16'd40462;
9'd442:value_o <=    16'd40723;
9'd443:value_o <=    16'd40988;
9'd444:value_o <=    16'd41256;
9'd445:value_o <=    16'd41528;
9'd446:value_o <=    16'd41803;
9'd447:value_o <=    16'd42082;
9'd448:value_o <=    16'd42365;
9'd449:value_o <=    16'd42651;
9'd450:value_o <=    16'd42940;
9'd451:value_o <=    16'd43233;
9'd452:value_o <=    16'd43530;
9'd453:value_o <=    16'd43829;
9'd454:value_o <=    16'd44132;
9'd455:value_o <=    16'd44438;
9'd456:value_o <=    16'd44748;
9'd457:value_o <=    16'd45060;
9'd458:value_o <=    16'd45375;
9'd459:value_o <=    16'd45694;
9'd460:value_o <=    16'd46015;
9'd461:value_o <=    16'd46340;
9'd462:value_o <=    16'd46667;
9'd463:value_o <=    16'd46997;
9'd464:value_o <=    16'd47330;
9'd465:value_o <=    16'd47666;
9'd466:value_o <=    16'd48004;
9'd467:value_o <=    16'd48346;
9'd468:value_o <=    16'd48689;
9'd469:value_o <=    16'd49035;
9'd470:value_o <=    16'd49384;
9'd471:value_o <=    16'd49735;
9'd472:value_o <=    16'd50089;
9'd473:value_o <=    16'd50444;
9'd474:value_o <=    16'd50802;
9'd475:value_o <=    16'd51163;
9'd476:value_o <=    16'd51525;
9'd477:value_o <=    16'd51890;
9'd478:value_o <=    16'd52256;
9'd479:value_o <=    16'd52625;
9'd480:value_o <=    16'd52995;
9'd481:value_o <=    16'd53368;
9'd482:value_o <=    16'd53742;
9'd483:value_o <=    16'd54118;
9'd484:value_o <=    16'd54496;
9'd485:value_o <=    16'd54875;
9'd486:value_o <=    16'd55256;
9'd487:value_o <=    16'd55639;
9'd488:value_o <=    16'd56023;
9'd489:value_o <=    16'd56409;
9'd490:value_o <=    16'd56795;
9'd491:value_o <=    16'd57184;
9'd492:value_o <=    16'd57573;
9'd493:value_o <=    16'd57964;
9'd494:value_o <=    16'd58356;
9'd495:value_o <=    16'd58748;
9'd496:value_o <=    16'd59142;
9'd497:value_o <=    16'd59537;
9'd498:value_o <=    16'd59933;
9'd499:value_o <=    16'd60330;
9'd500:value_o <=    16'd60727;
9'd501:value_o <=    16'd61125;
9'd502:value_o <=    16'd61524;
9'd503:value_o <=    16'd61923;
9'd504:value_o <=    16'd62323;
9'd505:value_o <=    16'd62724;
9'd506:value_o <=    16'd63124;
9'd507:value_o <=    16'd63526;
9'd508:value_o <=    16'd63927;
9'd509:value_o <=    16'd64329;
9'd510:value_o <=    16'd64731;
9'd511:value_o <=    16'd65133;
           default:   value_o <= 16'd0;
      endcase
 end    
endmodule  